.title KiCad schematic
U2 GND +3V3 Net-_C1-Pad1_ NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 GND NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 NC_19 NC_20 TOUCH_0 NC_21 NC_22 NC_23 NC_24 LED_DO LED_W NC_25 LED_B RX TX LED_G LED_R GND GND ESP32-WROOM
J1 B GND Conn_Coaxial_Power
U1 GND +3V3 B AMS1117-3.3
R1 +3V3 Net-_C1-Pad1_ 10k
C2 GND +3V3 10uF
C3 GND +3V3 100nF
SW1 Net-_C1-Pad1_ GND SW_Push
SW2 TOUCH_0 GND SW_Push
C1 Net-_C1-Pad1_ GND 100nF
Q1 LED_R B GND IRLB8721PBF
Q2 LED_G B GND IRLB8721PBF
Q3 LED_B B GND IRLB8721PBF
Q4 LED_W B GND IRLB8721PBF
TP1 LED_R TestPoint
TP3 LED_G TestPoint
TP5 LED_B TestPoint
TP7 LED_W TestPoint
TP2 B TestPoint
TP4 B TestPoint
TP6 B TestPoint
TP8 B TestPoint
J2 B B B B B Conn_01x05
Q5 LED_DO B GND IRLB8721PBF
TP9 LED_DO TestPoint
JP1 B DO LED_DO SolderJumper_3_Open
TP10 DO TestPoint
J3 B DO GND Conn_01x03
J4 +3V3 TX RX GND Conn_01x04
.end
